`timescale 1ns / 1ps

module Shift_ALU(clk,
           ALU_OP,
           A,
           B,
           Shift_Carry_Out,
           CF,
           VF,
           NZCV,
           F);
endmodule